`timescale 1ns / 1ps

////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer:
//
// Create Date:   11:03:41 05/02/2023
// Design Name:   stopwatch
// Module Name:   C:/Users/Student/Desktop/152alab10am/lab3/stopwatch_tb.v
// Project Name:  lab3
// Target Device:  
// Tool versions:  
// Description: 
//
// Verilog Test Fixture created by ISE for module: stopwatch
//
// Dependencies:
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
////////////////////////////////////////////////////////////////////////////////

module stopwatch_tb;

//	// Outputs
//	wire ;
//
//	// Instantiate the Unit Under Test (UUT)
//	stopwatch uut (
//		.()
//	);
//
//	initial begin
//		// Initialize Inputs
//
//		// Wait 100 ns for global reset to finish
//		#100;
//        
//		// Add stimulus here
//
//	end
      
endmodule

