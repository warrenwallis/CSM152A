module counter (
    input clk,
    input adj,
    input sel,
    input pse,
    input rst,
    output reg [3:0] sec_one,
    output reg [3:0] sec_ten,
    output reg [3:0] min_one,
    output reg [3:0] min_ten
);
    initial sec_one = 4'b0000;
    initial sec_ten = 4'b0000;
    initial min_one = 4'b0000;
    initial min_ten = 4'b0000;
    
    always @ (posedge clk or posedge rst) begin
             
        if (rst == 1'b1) begin // reset is pressed
            sec_one = 4'b0000;
            sec_ten = 4'b0000;
            min_one = 4'b0000;
            min_ten = 4'b0000;
        end
        
        else begin
            if (pse == 1'b0) begin
                // ADJ is LOW, stopwatch behaves normally
                if (adj == 1'b0) begin
                    if (sec_one < 10) begin
                        sec_one = sec_one + 1'b1;
                    end
                    else begin
                        sec_one = 4'b0000;
                        if (sec_ten < 6) begin
                            sec_ten = sec_ten + 1'b1;
                        end
                        else begin
                            sec_ten = 4'b0000;
                            if(min_one < 10) begin
                                min_one = min_one + 1'b1;
                            end
                            else begin
                                min_one = 4'b0000;
                                if (min_ten < 6) begin
                                    min_ten = min_ten + 1'b1;
                                end
                                else begin
                                    min_ten = 4'b0000;
                                end
                            end
                        end
                    end
                end
                // ADJ is HIGH, only increase selected digit
                else begin
                    if (sel == 1'b0) begin
                        if (min_one < 10) begin
                            min_one = min_one + 1'b1;
                        end
                        else begin
                            min_one = 4'b0000;
                            if (min_ten < 6) begin
                                min_ten = min_ten + 1'b1;
                            end
                            else begin
                                min_ten = 4'b0000;
                            end
                        end
                    end
                    else begin
                        // sec selected
                        if (sec_one < 10) begin
                            sec_one = sec_one + 1'b1;
                        end
                        else begin
                            sec_one = 4'b0000;
                            if (sec_ten < 6) begin
                                sec_ten = sec_ten + 1'b1;
                            end
                            else begin
                                sec_ten = 4'b0000;
                            end
                        end
                    end
                end
            end
        end
    end
    
endmodule
