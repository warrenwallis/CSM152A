module Stopwatch ();

endmodule