module display (
  //outputs
  sec, min,
  
  //inputs
  time
);
  
  output integer sec;
  output integer min;
  
  
  input time;
  
  always @ (posedge clk) begin
    
  end
  
endmodule
